
module SystemClk (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
